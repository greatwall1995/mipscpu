`include "defines.v"

module ex(  
  
    input wire             rst,  
      
    // ����׶��͵�ִ�н׶ε���Ϣ  
    input wire[`AluOpBus]         aluop_i,  
    input wire[`AluSelBus]        alusel_i,  
    input wire[`RegBus]           reg1_i,  
    input wire[`RegBus]           reg2_i,  
    input wire[`RegAddrBus]       wd_i,  
    input wire                    wreg_i,  
  
    // ִ�еĽ��  
    output reg[`RegAddrBus]       wd_o,  
    output reg                    wreg_o,  
    output reg[`RegBus]         wdata_o  
      
);  

	// �����߼�����Ľ��  
	reg[`RegBus] logicout;  
  
/****************************************************************** 
**  ��һ�Σ�����aluop_iָʾ�����������ͽ������㣬�˴�ֻ���߼��������� ** 
*******************************************************************/  

	always @ (*) begin  
		if(rst == `RstEnable) begin  
			logicout <= `ZeroWord;  
		end else begin  
			case (aluop_i)
				`EXE_AND_OP: begin
					logicout <= reg1_i & reg2_i;
				end
				`EXE_OR_OP: begin  
					logicout <= reg1_i | reg2_i;  
				end  
				`EXE_XOR_OP: begin
					logicout <= reg1_i ^ reg2_i;
				end
				default:    begin  
					logicout <= `ZeroWord;  
				end  
			endcase  
		end    //if  
	end      //always  
  
/**************************************************************** 
**  �ڶ��Σ�����alusel_iָʾ���������ͣ�ѡ��һ����������Ϊ���ս�� ** 
**         �˴�ֻ���߼�������                                 ** 
*****************************************************************/  
  
	always @ (*) begin  
		wd_o   <= wd_i;             // wd_o����wd_i��Ҫд��Ŀ�ļĴ�����ַ  
		wreg_o <= wreg_i;           // wreg_o����wreg_i����ʾ�Ƿ�ҪдĿ�ļĴ���  
		case ( alusel_i )   
			`EXE_RES_LOGIC: begin  
				wdata_o <= logicout;    // wdata_o�д��������
			end  
			default: begin  
				wdata_o <= `ZeroWord;  
			end  
		endcase  
	end
endmodule  