`include "defines.v"

module mem(  
  
    input wire           rst,  
      
    // ����ִ�н׶ε���Ϣ      
    input wire[`RegAddrBus]      wd_i,  
    input wire                   wreg_i,  
    input wire[`RegBus]      wdata_i,  
      
    // �ô�׶εĽ��  
    output reg[`RegAddrBus]      wd_o,  
    output reg                   wreg_o,  
    output reg[`RegBus]      wdata_o  
      
);  
  
    always @ (*) begin  
      if(rst == `RstEnable) begin  
        wd_o    <= `NOPRegAddr;  
        wreg_o  <= `WriteDisable;  
        wdata_o <= `ZeroWord;  
      end else begin  
        wd_o    <= wd_i;  
        wreg_o  <= wreg_i;  
        wdata_o <= wdata_i;  
      end      
    end        
  
endmodule  